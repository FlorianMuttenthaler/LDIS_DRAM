-------------------------------------------------------------------------------
--
-- KDF
--
-------------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--
-------------------------------------------------------------------------------
--
entity memory is

	-- is the generic value of the entity.
	-- are the inputs of entity.
	-- are the outputs of the entity.

	generic(
			
		);
		
	port (
		
	);

end memory;
--
-------------------------------------------------------------------------------
--
architecture beh of memory is

	
begin
	
--	slowclk: entity work.slowclk
--		port map(
--			R2 => R2,
--			R1 => R1,
--			X => X,			
--			clk_slow => clk_slow
--		);
	
end beh;
--
-------------------------------------------------------------------------------