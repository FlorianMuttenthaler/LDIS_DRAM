-------------------------------------------------------------------------------
--
-- 7-segment display package
--
-------------------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--
-------------------------------------------------------------------------------
--
package memory_pkg is

	component memory is

	-- is the generic value of the entity.
	-- are the inputs of entity.
	--  are the output of the entity.

	generic(

	);
		
	port (	

	);
	
	end component memory;
	
end memory_pkg;

